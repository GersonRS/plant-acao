1
7
vk
1
16
victor
1
10
Gerson
1
15
Gerson
1
31
Gerson
1
33
victor
1
0
Nenhum
1
11
Gerson
1
0
Nenhum
1
0
Nenhum